pb_top (
  input logic pclk,
  input logic preset_n,
  
  // Master inputs
  input logic [1:0] add_i,              // 2'b00 - NOP, 2'b01 - READ, 2'b11 - WRITE
  input logic [31:0] external_wdata_i,  // External write data
  
  // Outputs
  output logic ready_o,       // Slave ready signal
  output logic [31:0] rdata_o // Read data from slave
);

  // Declare and instantiate the APB interface
  apb_interface apb_intf (
    .pclk(pclk),
    .preset_n(preset_n)
  );

  // Instantiate the APB master using the master modport
  apb_master u_master (
    .add_i(add_i),
    .external_wdata_i(external_wdata_i),
    .apb_intf(apb_intf.master)  // Use the master modport
  );

  // Instantiate the APB slave using the slave modport
  apb_slave u_slave (
    .apb_intf(apb_intf.slave)   // Use the slave modport
  );

  // Connect outputs to the appropriate signals in the interface
  assign ready_o = apb_intf.pready;
  assign rdata_o = apb_intf.prdata;

endmodule

